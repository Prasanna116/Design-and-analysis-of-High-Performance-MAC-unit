module Wallace_Mult16(
input [15:0]a,
input [15:0]b,
output [31:0] out);

wire p[15:0][15:0];
wire cout;
wire [250:0]s,c;
wire [59:0] dot,ss,cc;
wire [31:0]z1,z2;

genvar i,j;
generate
for(i=0;i<16;i=i+1)begin :pp1
  for(j=0;j<16;j=j+1) begin:pp2
    assign p[j][i]=a[j] & b[i] ;
  end
end
endgenerate


// LEVEL 1 


assign dot[0] = p[0][0];
half_adder g1(p[1][0],p[0][1],ss[0],cc[0]);
full_adder g2(p[2][0],p[1][1],p[0][2],s[0],c[0]);
full_adder g3(p[3][0],p[2][1],p[1][2],s[1],c[1]);
full_adder g4(p[4][0],p[3][1],p[2][2],s[2],c[2]);
full_adder g5(p[5][0],p[4][1],p[3][2],s[3],c[3]);
full_adder g6(p[6][0],p[5][1],p[4][2],s[4],c[4]);
full_adder g7(p[7][0],p[6][1],p[5][2],s[5],c[5]);
full_adder g8(p[8][0],p[7][1],p[6][2],s[6],c[6]);
full_adder g9(p[9][0],p[8][1],p[7][2],s[7],c[7]);
full_adder g10(p[10][0],p[9][1],p[8][2],s[8],c[8]);
full_adder g11(p[11][0],p[10][1],p[9][2],s[9],c[9]);
full_adder g12(p[12][0],p[11][1],p[10][2],s[10],c[10]);
full_adder g13(p[13][0],p[12][1],p[11][2],s[11],c[11]);
full_adder g14(p[14][0],p[13][1],p[12][2],s[12],c[12]);
full_adder g15(p[15][0],p[14][1],p[13][2],s[13],c[13]);
half_adder g16(p[15][1],p[14][2],ss[1],cc[1]);
assign dot[1] = p[2][15];

assign dot[2] = p[3][0];
half_adder g17(p[1][3],p[0][4],ss[2],cc[2]);
full_adder g18(p[2][3],p[1][4],p[0][5],s[14],c[14]);
full_adder g19(p[3][3],p[2][4],p[1][5],s[15],c[15]);
full_adder g20(p[4][3],p[3][4],p[2][5],s[16],c[16]);
full_adder g21(p[5][3],p[4][4],p[3][5],s[17],c[17]);
full_adder g22(p[6][3],p[5][4],p[4][5],s[18],c[18]);
full_adder g23(p[7][3],p[6][4],p[5][5],s[19],c[19]);
full_adder g24(p[8][3],p[7][4],p[6][5],s[20],c[20]);
full_adder g25(p[9][3],p[8][4],p[7][5],s[21],c[21]);
full_adder g26(p[10][3],p[9][4],p[8][5],s[22],c[22]);
full_adder g27(p[11][3],p[10][4],p[9][5],s[23],c[23]);
full_adder g28(p[12][3],p[11][4],p[10][5],s[24],c[24]);
full_adder g29(p[13][3],p[12][4],p[11][5],s[25],c[25]);
full_adder g30(p[14][3],p[13][4],p[12][5],s[26],c[26]);
full_adder g31(p[15][3],p[14][4],p[13][5],s[27],c[27]);
half_adder g32(p[15][4],p[14][5],ss[3],cc[3]);
assign dot[3]=p[15][5];

assign dot[4] = p[0][6];
half_adder g33(p[1][6],p[0][7],ss[4],cc[4]);
full_adder g34(p[2][6],p[1][7],p[0][8],s[28],c[28]);
full_adder g35(p[3][6],p[2][7],p[1][8],s[29],c[29]);
full_adder g36(p[4][6],p[3][7],p[2][8],s[30],c[30]);
full_adder g37(p[5][6],p[4][7],p[3][8],s[31],c[31]);
full_adder g38(p[6][6],p[5][7],p[4][8],s[32],c[32]);
full_adder g39(p[7][6],p[6][7],p[5][8],s[33],c[33]);
full_adder g40(p[8][6],p[7][7],p[6][8],s[34],c[34]);
full_adder g41(p[9][6],p[8][7],p[7][8],s[35],c[35]);
full_adder g42(p[10][6],p[9][7],p[8][8],s[36],c[36]);
full_adder g43(p[11][6],p[10][7],p[9][8],s[37],c[37]);
full_adder g44(p[12][6],p[11][7],p[10][8],s[38],c[38]);
full_adder g45(p[13][6],p[12][7],p[11][8],s[39],c[39]);
full_adder g46(p[14][6],p[13][7],p[12][8],s[40],c[40]);
full_adder g47(p[15][6],p[14][7],p[13][8],s[41],c[41]);
half_adder g48(p[15][7],p[14][8],ss[5],cc[5]);
assign dot[5] = p[15][8];

assign dot[6] = p[0][9];
half_adder g49(p[1][9],p[0][10],ss[6],cc[6]);
full_adder g50(p[2][9],p[1][10],p[0][11],s[42],c[42]);
full_adder g51(p[3][9],p[2][10],p[1][11],s[43],c[43]);
full_adder g52(p[4][9],p[3][10],p[2][11],s[44],c[44]);
full_adder g53(p[5][9],p[4][10],p[3][11],s[45],c[45]);
full_adder g54(p[6][9],p[5][10],p[4][11],s[46],c[46]);
full_adder g55(p[7][9],p[6][10],p[5][11],s[47],c[47]);
full_adder g56(p[8][9],p[7][10],p[6][11],s[48],c[48]);
full_adder g57(p[9][9],p[8][10],p[7][11],s[49],c[49]);
full_adder g58(p[10][9],p[9][10],p[8][11],s[50],c[50]);
full_adder g59(p[11][9],p[10][10],p[9][11],s[51],c[51]);
full_adder g60(p[12][9],p[11][10],p[10][11],s[52],c[52]);
full_adder g61(p[13][9],p[12][10],p[11][11],s[53],c[53]);
full_adder g62(p[14][9],p[13][10],p[12][11],s[54],c[54]);
full_adder g63(p[15][9],p[14][10],p[13][11],s[55],c[55]);
half_adder g64(p[15][10],p[14][11],ss[7],cc[7]);
assign dot[7] = p[15][11];

assign dot[8] = p[0][12];
half_adder g65(p[1][12],p[0][13],ss[8],cc[8]);
full_adder g66(p[2][12],p[1][13],p[0][14],s[56],c[56]);
full_adder g67(p[3][12],p[2][13],p[1][14],s[57],c[57]);
full_adder g68(p[4][12],p[3][13],p[2][14],s[58],c[58]);
full_adder g69(p[5][12],p[4][13],p[3][14],s[59],c[59]);
full_adder g70(p[6][12],p[5][13],p[4][14],s[60],c[60]);
full_adder g71(p[7][12],p[6][13],p[5][14],s[61],c[61]);
full_adder g72(p[8][12],p[7][13],p[6][14],s[62],c[62]);
full_adder g73(p[9][12],p[8][13],p[7][14],s[63],c[63]);
full_adder g74(p[10][12],p[9][13],p[8][14],s[64],c[64]);
full_adder g75(p[11][12],p[10][13],p[9][14],s[65],c[65]);
full_adder g76(p[12][12],p[11][13],p[10][14],s[66],c[66]);
full_adder g77(p[13][12],p[12][13],p[11][14],s[67],c[67]);
full_adder g78(p[14][12],p[13][13],p[12][14],s[68],c[68]);
full_adder g79(p[15][12],p[14][13],p[13][14],s[69],c[69]);
half_adder g80(p[15][13],p[14][14],ss[9],cc[9]);
assign dot[9] = p[15][14];

assign dot[10] = p[0][15];
assign dot[11] = p[1][15];
assign dot[12] = p[2][15];
assign dot[13] = p[3][15];
assign dot[14] = p[4][15];
assign dot[15] = p[5][15];
assign dot[16] = p[6][15];
assign dot[17] = p[7][15];
assign dot[18] = p[8][15];
assign dot[19] = p[9][15];
assign dot[20] = p[10][15];
assign dot[21] = p[11][15];
assign dot[22] = p[12][15];
assign dot[23] = p[13][15];
assign dot[24] = p[14][15];
assign dot[25] = p[15][15];

//LEVEL 2

assign dot[26] = dot[0];
assign dot[27] = ss[0];

half_adder g81(s[0], cc[0], ss[10], cc[10]);
full_adder g82(s[1], c[0], dot[2], s[70], c[70]);
full_adder g83(s[2], c[1], ss[2], s[71], c[71]);
full_adder g84(s[3], c[2], s[14], s[72], c[72]);
full_adder g85(s[4], c[3], s[15], s[73], c[73]);
full_adder g86(s[5], c[4], s[16], s[74], c[74]);
full_adder g87(s[6], c[5], s[17], s[75], c[75]);
full_adder g88(s[7], c[6], s[18], s[76], c[76]);
full_adder g89(s[8], c[7], s[19], s[77], c[77]);
full_adder g90(s[9], c[8], s[20], s[78], c[78]);
full_adder g91(s[10], c[9], s[21], s[79], c[79]);
full_adder g92(s[11], c[10], s[23], s[80], c[80]);
full_adder g93(s[12], c[11], s[24], s[81], c[81]);
full_adder g94(s[13], c[12], s[25], s[82], c[82]);
full_adder g95(ss[1], c[13], s[26], s[83], c[83]);
full_adder g96(dot[1], cc[1], s[27], s[84], c[84]);
assign dot[28] = s[28];
assign dot[29] = ss[3];
assign dot[30] = dot[3];

assign dot[31] = cc[2];
half_adder g97(c[14], dot[4], ss[11], cc[11]);
half_adder g98(c[15], ss[4], ss[12], cc[12]);
full_adder g99(c[16], s[28], cc[4], s[85], c[85]);
full_adder g100(c[17], s[29], c[28], s[86], c[86]);
full_adder g101(c[18], s[30], c[29], s[87], c[87]);
full_adder g102(c[19], s[31], c[30], s[88], c[88]);
full_adder g103(c[20], s[32], c[31], s[89], c[89]);
full_adder g104(c[21], s[33], c[32], s[90], c[90]);
full_adder g105(c[22], s[34], c[33], s[91], c[91]);
full_adder g106(c[23], s[35], c[34], s[92], c[92]);
full_adder g107(c[24], s[36], c[35], s[93], c[93]);
full_adder g108(c[25], s[37], c[36], s[94], c[94]);
full_adder g109(c[26], s[38], c[37], s[95], c[95]);
full_adder g110(c[27], s[39], c[38], s[96], c[96]);
full_adder g111(cc[3], s[40], c[39], s[97], c[97]);
half_adder g112(s[41], c[40], ss[13], cc[13]);
half_adder g113(ss[5], c[41], ss[14], cc[14]);
half_adder g114(dot[5], cc[5], ss[15], cc[15]);

assign dot[32] = dot[6];
assign dot[33] = ss[6];
half_adder g115(s[42], cc[6], ss[16], cc[16]);
full_adder g116(s[43], c[42], dot[8], s[98], c[98]);
full_adder g117(s[44], c[43], ss[8], s[99], c[99]);
full_adder g118(s[45], c[44], s[56], s[100], c[100]);
full_adder g119(s[46], c[45], s[57], s[101], c[101]);
full_adder g120(s[47], c[46], s[58], s[102], c[102]);
full_adder g121(s[48], c[47], s[59], s[103], c[103]);
full_adder g122(s[49], c[48], s[60], s[104], c[104]);
full_adder g123(s[50], c[49], s[61], s[105], c[105]);
full_adder g124(s[51], c[50], s[62], s[106], c[106]);
full_adder g125(s[52], c[51], s[63], s[107], c[107]);
full_adder g126(s[53], c[52], s[64], s[108], c[108]);
full_adder g127(s[54], c[53], s[65], s[109], c[109]);
full_adder g128(s[55], c[54], s[66], s[110], c[110]);
full_adder g129(ss[7], c[55], s[67], s[111], c[111]);
full_adder g130(dot[7], cc[7], s[68], s[112], c[112]);
assign dot[34] = s[69];
assign dot[35] = ss[9];
assign dot[36] = dot[9];

//last two rows of dots will carry over a few times, keep track of them

//LEVEL 3
//dot[26], dot[27]
assign dot[37] = ss[10];
half_adder g131(s[70], cc[10], ss[17], cc[17]);
half_adder g132(s[71], c[70], ss[18], cc[18]);
full_adder g133(s[72], c[71], dot[31], s[113], c[113]);
full_adder g134(s[73], c[72], ss[11], s[114], c[114]);
full_adder g135(s[74], c[73], ss[12], s[115], c[115]);
full_adder g136(s[75], c[74], s[85], s[116], c[116]);
full_adder g137(s[76], c[75], s[86], s[117], c[117]);
full_adder g138(s[77], c[76], s[87], s[118], c[118]);
full_adder g139(s[78], c[77], s[88], s[119], c[119]);
full_adder g140(s[79], c[78], s[89], s[120], c[120]);
full_adder g141(s[80], c[79], s[90], s[121], c[121]);
full_adder g142(s[81], c[80], s[91], s[122], c[122]);
full_adder g143(s[82], c[81], s[92], s[123], c[123]);
full_adder g144(s[83], c[82], s[93], s[124], c[124]);
full_adder g145(s[84], c[83], s[94], s[125], c[125]);
full_adder g146(dot[28], c[84], s[95], s[126], c[126]);
half_adder g147(dot[29], s[96], ss[19], cc[19]);
half_adder g148(dot[30], s[97], ss[20], cc[20]);
assign dot[38] = ss[13];
assign dot[39] = ss[14];
assign dot[40] = ss[15];

assign dot[41] = cc[11];
assign dot[42] = cc[12];
half_adder g149(c[85], dot[32], ss[21], cc[21]);
half_adder g150(c[86], c[86], ss[22], cc[22]);
half_adder g151(c[87], ss[16], ss[23], cc[23]);
full_adder g152(c[88], s[98], cc[16], s[127], c[127]);
full_adder g153(c[89], s[99], c[98], s[128], c[128]);
full_adder g154(c[90], s[100], c[99], s[129], c[129]);
full_adder g155(c[91], s[101], c[100], s[130], c[130]);
full_adder g156(c[92], s[102], c[101], s[131], c[131]);
full_adder g157(c[93], s[103], c[102], s[132], c[132]);
full_adder g158(c[94], s[104], c[103], s[133], c[133]);
full_adder g159(c[95], s[105], c[104], s[134], c[134]);
full_adder g160(c[96], s[106], c[105], s[135], c[135]);
full_adder g161(c[97], s[107], c[106], s[136], c[136]);
full_adder g162(cc[13], s[108], c[107], s[137], c[137]);
full_adder g163(cc[14], s[109], c[108], s[138], c[138]);
full_adder g164(cc[15], s[110], c[109], s[139], c[139]);
half_adder g165(s[111], c[110], ss[24], cc[24]);
half_adder g166(s[112], c[111], ss[25], cc[25]);
half_adder g167(dot[34], c[112], ss[26], cc[26]);
assign dot[43] = dot[35];
assign dot[44] = dot[36];

/***************/

// LEVEL 4 
//dot[26], [27], [37]

assign dot[45] = ss[17];
half_adder g168(ss[18], cc[17], ss[27], cc[27]);
half_adder g169(s[113], cc[18], ss[28], cc[28]);
half_adder g170(s[114], c[113], ss[29], cc[29]);
full_adder g171(s[115], c[114], dot[41], s[140], c[140]);
full_adder g172(s[116], c[115], dot[42], s[141], c[141]);
full_adder g173(s[117], c[116], ss[21], s[142], c[142]);
full_adder g174(s[118], c[117], ss[22], s[143], c[143]);
full_adder g175(s[119], c[118], ss[23], s[144], c[144]);
full_adder g176(s[120], c[119], s[127], s[145], c[145]);
full_adder g177(s[121], c[120], s[128], s[146], c[146]);
full_adder g178(s[122], c[121], s[129], s[147], c[147]);
full_adder g179(s[123], c[122], s[130], s[148], c[148]);
full_adder g180(s[124], c[123], s[131], s[149], c[149]);
full_adder g181(s[125], c[124], s[132], s[150], c[150]);
full_adder g182(s[126], c[125], s[133], s[151], c[151]);
full_adder g183(ss[19], c[126], s[134], s[152], c[152]);
full_adder g184(ss[20], cc[19], s[135], s[153], c[153]);
full_adder g185(dot[38], cc[20], s[136], s[154], c[154]);
half_adder g186(dot[39], s[137], ss[30], cc[30]);
half_adder g187(dot[40], s[138], ss[31], cc[31]);
assign dot[46] = s[139];
assign dot[47] = ss[24];
assign dot[48] = ss[25];
assign dot[49] = ss[26];
//dot[43]

assign dot[50] = cc[21];
assign dot[51] = cc[22];
assign dot[52] = cc[23];
assign dot[53] = c[127];

half_adder g188(c[128], cc[8], ss[32], cc[32]); //check first for errors
full_adder g189(c[129], c[56], dot[10], s[155], c[155]);
full_adder g190(c[130], c[57], dot[11], s[156], c[156]);
full_adder g191(c[131], c[58], dot[12], s[157], c[157]);
full_adder g192(c[132], c[59], dot[13], s[158], c[158]);
full_adder g193(c[133], c[60], dot[14], s[159], c[159]);
full_adder g194(c[134], c[61], dot[15], s[160], c[160]);
full_adder g195(c[135], c[62], dot[16], s[161], c[161]);
full_adder g196(c[136], c[63], dot[17], s[162], c[162]);
full_adder g197(c[137], c[64], dot[18], s[163], c[163]);
full_adder g198(c[138], c[65], dot[19], s[164], c[164]);
full_adder g199(c[139], c[66], dot[20], s[165], c[165]);
full_adder g200(cc[24], c[67], dot[21], s[166], c[166]);
full_adder g201(cc[25], c[68], dot[22], s[167], c[167]);
full_adder g202(cc[26], c[69], dot[23], s[168], c[168]);
full_adder g203(dot[36], cc[9], dot[24], s[169], c[169]);
assign dot[54] = dot[25];

/**************/
// LEVEL 5
//dot[26], [27], [37], [45]

assign dot[55] = ss[27];
half_adder g204(ss[28], cc[27], ss[33], cc[33]);
half_adder g205(ss[29], cc[28], ss[34], cc[34]);
half_adder g206(s[140], cc[29], ss[35], cc[35]);
half_adder g207(s[141], c[140], ss[36], cc[36]);
half_adder g208(s[142], c[141], ss[37], cc[37]);
full_adder g209(s[143], c[142], dot[50], s[170], c[170]);
full_adder g210(s[144], c[143], dot[51], s[171], c[171]);
full_adder g211(s[145], c[144], dot[52], s[172], c[172]);
full_adder g212(s[146], c[145], dot[53], s[173], c[173]);
full_adder g213(s[147], c[146], ss[32], s[174], c[174]);
full_adder g214(s[148], c[147], s[155], s[175], c[175]);
full_adder g215(s[149], c[148], s[156], s[176], c[176]);
full_adder g216(s[150], c[149], s[157], s[177], c[177]);
full_adder g217(s[151], c[150], s[158], s[178], c[178]);
full_adder g218(s[152], c[151], s[159], s[179], c[179]);
full_adder g219(s[153], c[152], s[160], s[180], c[180]);
full_adder g220(s[154], c[153], s[161], s[181], c[181]);
full_adder g221(ss[30], c[154], s[162], s[182], c[182]);
full_adder g222(ss[31], cc[30], s[163], s[183], c[183]);
full_adder g223(dot[46], cc[31], s[164], s[184], c[184]);
half_adder g224(dot[47], s[165], ss[38], cc[38]);
half_adder g225(dot[48], s[166], ss[39], cc[39]);
half_adder g226(dot[49], s[167], ss[40], cc[40]);
half_adder g227(dot[43], s[168], ss[41], cc[41]);
assign dot[56] = s[169];

/*************/
// level 6

assign dot[57] = ss[33];
half_adder g228(ss[34], cc[33], ss[42], cc[42]);
half_adder g229(ss[35], cc[34], ss[43], cc[43]);
half_adder g230(ss[36], cc[35], ss[44], cc[44]);
half_adder g231(ss[37], cc[36], ss[45], cc[45]);
half_adder g232(s[170], cc[37], ss[46], cc[46]);
half_adder g233(s[171], c[170], ss[47], cc[47]);
half_adder g234(s[172], c[171], ss[48], cc[48]);
half_adder g235(s[173], c[172], ss[49], cc[49]);
half_adder g236(s[174], c[173], ss[50], cc[50]);
full_adder g237(s[175], c[174], cc[32], s[185], c[185]);
full_adder g238(s[176], c[175], c[155], s[186], c[186]);
full_adder g239(s[177], c[176], c[156], s[187], c[187]);
full_adder g240(s[178], c[177], c[157], s[188], c[188]);
full_adder g241(s[179], c[178], c[158], s[189], c[189]);
full_adder g242(s[180], c[179], c[159], s[190], c[190]);
full_adder g243(s[181], c[180], c[160], s[191], c[191]);
full_adder g244(s[182], c[181], c[161], s[192], c[192]);
full_adder g245(s[183], c[182], c[162], s[193], c[193]);
full_adder g246(s[184], c[183], c[163], s[194], c[194]);
full_adder g247(ss[38], c[184], c[164], s[195], c[195]);
full_adder g248(ss[39], cc[38], c[165], s[196], c[196]);
full_adder g249(ss[40], cc[39], c[166], s[197], c[197]);
full_adder g250(ss[41], cc[40], c[167], s[198], c[198]);
full_adder g251(dot[56], cc[41], c[168], s[199], c[199]);
half_adder g252(dot[54], c[169], ss[51], cc[51]);

/*************/
//LEVEL 7

assign z1[0] = dot[26];
assign z1[1] = dot[27];
assign z1[2] = dot[37];
assign z1[3] = dot[45];
assign z1[4] = dot[55];
assign z1[5] = dot[57];
assign z1[6] = ss[42];
assign z1[7] = ss[43];
assign z1[8] = ss[44];
assign z1[9] = ss[45];
assign z1[10] = ss[46];
assign z1[11] = ss[47];
assign z1[12] = ss[48];
assign z1[13] = ss[49];
assign z1[14] = ss[50];
assign z1[15] = s[185];
assign z1[16] = s[186];
assign z1[17] = s[187];
assign z1[18] = s[188];
assign z1[19] = s[189];
assign z1[20] = s[190];
assign z1[21] = s[191];
assign z1[22] = s[192];
assign z1[23] = s[193];
assign z1[24] = s[194];
assign z1[25] = s[195];
assign z1[26] = s[196];
assign z1[27] = s[197];
assign z1[28] = s[198];
assign z1[29] = s[199];
assign z1[30] = ss[51];
assign z1[31] = 0;

assign z2[0] = 0;
assign z2[1] = 0;
assign z2[2] = 0;
assign z2[3] = 0;
assign z2[4] = 0;
assign z2[5] = 0;
assign z2[6] = 0;
assign z2[7] = cc[42];
assign z2[8] = cc[43];
assign z2[9] = cc[44];
assign z2[10] = cc[45];
assign z2[11] = cc[46];
assign z2[12] = cc[47];
assign z2[13] = cc[48];
assign z2[14] = cc[49];
assign z2[15] = cc[50];
assign z2[16] = c[185];
assign z2[17] = c[186];
assign z2[18] = c[187];
assign z2[19] = c[188];
assign z2[20] = c[189];
assign z2[21] = c[190];
assign z2[22] = c[191];
assign z2[23] = c[192];
assign z2[24] = c[193];
assign z2[25] = c[194];
assign z2[26] = c[195];
assign z2[27] = c[196];
assign z2[28] = c[197];
assign z2[29] = c[198];
assign z2[30] = c[199];
assign z2[31] = cc[51];

assign out[0]=z1[0];
assign out[1]=z1[1];
assign out[2]=z1[2];
assign out[3]=z1[3];
assign out[4]=z1[4];
assign out[5]=z1[5];
assign out[6]=z1[6];

half_adder gg54(z1[7],z2[7],out[7],c[200]);
full_adder gg55(z1[8],z2[8],c[200],out[8],c[201]);
full_adder gg56(z1[9],z2[9],c[201],out[9],c[202]);
full_adder gg57(z1[10],z2[10],c[202],out[10],c[203]);
full_adder gg58(z1[11], z2[11], c[203], out[11], c[204]);
full_adder gg59(z1[12], z2[12], c[204], out[12], c[205]);
full_adder gg60(z1[13], z2[13], c[205], out[13], c[206]);
full_adder gg61(z1[14], z2[14], c[206], out[14], c[207]);
full_adder gg62(z1[15], z2[15], c[207], out[15], c[208]);
full_adder gg63(z1[16], z2[16], c[208], out[16], c[209]);
full_adder gg64(z1[17], z2[17], c[209], out[17], c[210]);
full_adder gg65(z1[18], z2[18], c[210], out[18], c[211]);
full_adder gg66(z1[19], z2[19], c[211], out[19], c[212]);
full_adder gg67(z1[20], z2[20], c[212], out[20], c[213]);
full_adder gg68(z1[21], z2[21], c[213], out[21], c[214]);
full_adder gg69(z1[22], z2[22], c[214], out[22], c[215]);
full_adder gg70(z1[23], z2[23], c[215], out[23], c[216]);
full_adder gg71(z1[24], z2[24], c[216], out[24], c[217]);
full_adder gg72(z1[25], z2[25], c[217], out[25], c[218]);
full_adder gg73(z1[26], z2[26], c[218], out[26], c[219]);
full_adder gg74(z1[27], z2[27], c[219], out[27], c[220]);
full_adder gg75(z1[28], z2[28], c[220], out[28], c[221]);
full_adder gg76(z1[29], z2[29], c[221], out[29], c[222]);
full_adder gg77(z1[30], z2[30], c[222], out[30], c[223]);
half_adder gg78(z2[31], c[223], out[31], c[224]);  // Final carry in = c[223]


//CarryLookAhead32_Adder ytt(z1[31:0],z2[31:0],0,out,cout);

endmodule

